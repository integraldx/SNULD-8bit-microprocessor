`timescale 1ns/1ps

module controller
(
    input [1:0] mode,
    input [1:0] opcode,
    output register_write,
    output memory_write,
    output pc_write,
    output memory_to_register,
    output alu_negation,
);
    

endmodule